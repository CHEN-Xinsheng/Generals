module Random_Boards_Library
#(parameter WORDS_CNT = 4096) (
    input wire [$clog2(WORDS_CNT) - 1: 0] address,
    output wire [3:0] h,
    output wire [3:0] v,
    output wire [1:0] piece_type
);

assign h            = init_boards[address][9:6];
assign v            = init_boards[address][5:2];
assign piece_type   = init_boards[address][1:0];

localparam [0:4095][9:0] init_boards = {
    10'b0001001110,
    10'b1000100011,
    10'b0001100100,
    10'b0110000000,
    10'b1000000000,
    10'b1001011000,
    10'b0111010100,
    10'b0100000000,
    10'b0011011100,
    10'b1001010000,
    10'b0010010000,
    10'b0000100100,
    10'b1001001100,
    10'b1000100100,
    10'b0010001001,
    10'b1001100001,
    10'b0001001001,
    10'b0111010001,
    10'b1000001001,
    10'b0010001101,
    10'b1000010101,
    10'b0011001001,
    10'b0111100001,
    10'b0100010101,
    10'b0110011001,
    10'b0010000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000011010,
    10'b0001000111,
    10'b0011010100,
    10'b0100000100,
    10'b1001010000,
    10'b1000000100,
    10'b0001010000,
    10'b0110100100,
    10'b0011000000,
    10'b0111000000,
    10'b0011001100,
    10'b0110010100,
    10'b0101011100,
    10'b0000100100,
    10'b0100011100,
    10'b0001001000,
    10'b0111100000,
    10'b1001011001,
    10'b0010001001,
    10'b0101010001,
    10'b0010011001,
    10'b0011001001,
    10'b1001100001,
    10'b0101000001,
    10'b0001100001,
    10'b0000010001,
    10'b1001001101,
    10'b1001001001,
    10'b0010001101,
    10'b0111010001,
    10'b0010100001,
    10'b0010011101,
    10'b0001100010,
    10'b0111000111,
    10'b0010000000,
    10'b0111011000,
    10'b0001000100,
    10'b0101001100,
    10'b0000010100,
    10'b0011010000,
    10'b0111011100,
    10'b1001011100,
    10'b0001011000,
    10'b1000000000,
    10'b1000100000,
    10'b1000000100,
    10'b0101011000,
    10'b1000011100,
    10'b0000011101,
    10'b1000001001,
    10'b0011000101,
    10'b0001010001,
    10'b0010011001,
    10'b0011001101,
    10'b0100011001,
    10'b0101010001,
    10'b0110100001,
    10'b0001001101,
    10'b0011011001,
    10'b1000010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000001011,
    10'b1001100000,
    10'b0110000100,
    10'b0000010000,
    10'b1001100100,
    10'b1001010000,
    10'b0000100000,
    10'b0110100000,
    10'b0101100100,
    10'b0110010100,
    10'b0100000000,
    10'b1000011100,
    10'b0111100100,
    10'b0100000100,
    10'b0001100101,
    10'b0111001001,
    10'b0011000001,
    10'b0100011001,
    10'b0111000101,
    10'b0000000001,
    10'b1000100001,
    10'b0011001101,
    10'b0000010101,
    10'b0100010101,
    10'b0111100001,
    10'b1000000101,
    10'b0101001101,
    10'b0100010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001100011,
    10'b0000100100,
    10'b1001011100,
    10'b1000001000,
    10'b0100001000,
    10'b0110000100,
    10'b0010100100,
    10'b1000011100,
    10'b0011001100,
    10'b1001001100,
    10'b0100100100,
    10'b1000000000,
    10'b1000001001,
    10'b0010011101,
    10'b0111010001,
    10'b0000000001,
    10'b0111100001,
    10'b0111001101,
    10'b0111000101,
    10'b1001010101,
    10'b0010001001,
    10'b0101000101,
    10'b0011000001,
    10'b1001000101,
    10'b0110001101,
    10'b0011010001,
    10'b0101001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001011111,
    10'b0010000100,
    10'b0111010100,
    10'b1000000000,
    10'b0001010000,
    10'b1001000100,
    10'b0000000000,
    10'b1001001000,
    10'b0011010000,
    10'b0110010100,
    10'b0101000100,
    10'b0110011100,
    10'b0000011000,
    10'b0101000000,
    10'b1000100000,
    10'b1000010100,
    10'b1000001101,
    10'b0010100001,
    10'b0111001001,
    10'b1001011101,
    10'b0000001001,
    10'b0010100101,
    10'b1000000101,
    10'b0101001101,
    10'b0000100001,
    10'b0101010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001100011,
    10'b0111000000,
    10'b0100011000,
    10'b0000011000,
    10'b0101001100,
    10'b1001011100,
    10'b1001010000,
    10'b1001100000,
    10'b0100000100,
    10'b0101010100,
    10'b0110011100,
    10'b0000001100,
    10'b0000100000,
    10'b0001011000,
    10'b0000000000,
    10'b0100001000,
    10'b0000000100,
    10'b1000011100,
    10'b1000011000,
    10'b1000000101,
    10'b0010100001,
    10'b0101000101,
    10'b0101011001,
    10'b0000010001,
    10'b0110000101,
    10'b0011010101,
    10'b0000100101,
    10'b0011010001,
    10'b0010010001,
    10'b1001011001,
    10'b1111111100,
    10'b0001000110,
    10'b1000100011,
    10'b0000001000,
    10'b0001010000,
    10'b0010100000,
    10'b0010011100,
    10'b0111000000,
    10'b0101011100,
    10'b0111100000,
    10'b1000000100,
    10'b1001010000,
    10'b0010010100,
    10'b0001011000,
    10'b0110001000,
    10'b0110100100,
    10'b0101000000,
    10'b0110010100,
    10'b0001001001,
    10'b0111100101,
    10'b0010001001,
    10'b0010100101,
    10'b0100011001,
    10'b0111011101,
    10'b0111011001,
    10'b0100010101,
    10'b1000011101,
    10'b0011100101,
    10'b0001100001,
    10'b0110001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000000111,
    10'b0001100100,
    10'b1001000000,
    10'b0001010000,
    10'b0101011100,
    10'b0100011000,
    10'b0011000000,
    10'b1000011000,
    10'b1000011100,
    10'b1000001000,
    10'b0100011100,
    10'b0100001100,
    10'b0000001000,
    10'b0001000000,
    10'b0000100101,
    10'b1001000001,
    10'b1001001001,
    10'b0111100101,
    10'b0011000101,
    10'b0011001101,
    10'b1000001101,
    10'b0100010101,
    10'b0100000101,
    10'b0100100101,
    10'b0001010101,
    10'b0110100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010100010,
    10'b1000001011,
    10'b0001001000,
    10'b0001000000,
    10'b1001100100,
    10'b0111000000,
    10'b1001001000,
    10'b0011001000,
    10'b0000011000,
    10'b0101100000,
    10'b1001000100,
    10'b0100100100,
    10'b0011001100,
    10'b0000100000,
    10'b0111000100,
    10'b0011000000,
    10'b0011100001,
    10'b0111001101,
    10'b0011011001,
    10'b1000000001,
    10'b0011010101,
    10'b0000001101,
    10'b0000000001,
    10'b0000100101,
    10'b0010100101,
    10'b1000001101,
    10'b0001100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001001110,
    10'b1000100011,
    10'b0100001100,
    10'b0001010000,
    10'b0111001100,
    10'b0010100100,
    10'b0010000100,
    10'b0011010100,
    10'b0111011100,
    10'b0011100000,
    10'b0110010000,
    10'b0101011100,
    10'b0000010001,
    10'b0111011101,
    10'b0000100101,
    10'b1001100101,
    10'b1000010001,
    10'b0111100101,
    10'b0100010001,
    10'b0000000101,
    10'b0100001001,
    10'b0010100001,
    10'b0011000001,
    10'b0110100101,
    10'b1001011001,
    10'b0101010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0011000111,
    10'b1000000100,
    10'b0110000000,
    10'b1000011000,
    10'b0011001100,
    10'b1000001100,
    10'b0111010000,
    10'b0110000100,
    10'b0110001000,
    10'b1001100000,
    10'b0000100100,
    10'b0101100000,
    10'b0010010100,
    10'b1001011101,
    10'b0100001001,
    10'b0111000001,
    10'b1001010101,
    10'b0110011001,
    10'b0111100101,
    10'b0100000101,
    10'b0000011101,
    10'b0000000001,
    10'b1001001001,
    10'b0111001101,
    10'b0011001001,
    10'b0001011101,
    10'b0010001001,
    10'b0001011001,
    10'b0110100101,
    10'b1000010001,
    10'b1111111100,
    10'b0111000110,
    10'b0001011111,
    10'b1000001100,
    10'b1001011000,
    10'b0010000000,
    10'b0100010000,
    10'b1000100100,
    10'b0011000100,
    10'b1000011000,
    10'b0010100100,
    10'b1001000100,
    10'b0000010000,
    10'b0011010000,
    10'b1001010000,
    10'b0000011000,
    10'b0001001100,
    10'b0111000001,
    10'b0001011001,
    10'b1001001001,
    10'b0100000001,
    10'b0010001101,
    10'b1001100101,
    10'b0001000101,
    10'b0000001001,
    10'b0100100101,
    10'b0111011001,
    10'b0100100001,
    10'b0101011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b0110100011,
    10'b1000001100,
    10'b0001011100,
    10'b0010011000,
    10'b0011100100,
    10'b0001100100,
    10'b0100000100,
    10'b0110001100,
    10'b1000010100,
    10'b0101010000,
    10'b0101011100,
    10'b1000001000,
    10'b0000000000,
    10'b0101001000,
    10'b0000000101,
    10'b0101100101,
    10'b0011001101,
    10'b0110100101,
    10'b0110001001,
    10'b0111000001,
    10'b0110000001,
    10'b0010010101,
    10'b1000011101,
    10'b0011000101,
    10'b0110000101,
    10'b0010010001,
    10'b0100100101,
    10'b0110010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0011000111,
    10'b0111010000,
    10'b0101000000,
    10'b1001100000,
    10'b1000000000,
    10'b1000001100,
    10'b0101000100,
    10'b1001010000,
    10'b0011010000,
    10'b0001001000,
    10'b0000010000,
    10'b0110011100,
    10'b0111100000,
    10'b1001001100,
    10'b0000011000,
    10'b1000000100,
    10'b0001100000,
    10'b0011001100,
    10'b0001000100,
    10'b0110001000,
    10'b1000100101,
    10'b0011001001,
    10'b0010010101,
    10'b0001000001,
    10'b1001010101,
    10'b0110100001,
    10'b0101001001,
    10'b0100100101,
    10'b0111011001,
    10'b0001011001,
    10'b0100100001,
    10'b0001001010,
    10'b1000100011,
    10'b0000001000,
    10'b1001011100,
    10'b0110100000,
    10'b1001000000,
    10'b0001011100,
    10'b0100000000,
    10'b1000011000,
    10'b0100011100,
    10'b0010001100,
    10'b0101001100,
    10'b0010100100,
    10'b0000000101,
    10'b1001100101,
    10'b0101000101,
    10'b0011010101,
    10'b0011001001,
    10'b0001001101,
    10'b0100001001,
    10'b0111001101,
    10'b1001011001,
    10'b0111100001,
    10'b0000100101,
    10'b0100010101,
    10'b0100100001,
    10'b0101100001,
    10'b0011010001,
    10'b0100100101,
    10'b0110011101,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001100011,
    10'b0100000000,
    10'b0100100100,
    10'b0110001000,
    10'b1001011100,
    10'b1001010000,
    10'b0111011100,
    10'b0110100000,
    10'b0110100100,
    10'b0101000000,
    10'b0000000100,
    10'b1000000101,
    10'b0001011101,
    10'b0010010101,
    10'b0000100101,
    10'b0100011101,
    10'b0101001001,
    10'b0111000001,
    10'b0110000101,
    10'b0010100101,
    10'b0111011001,
    10'b0101001101,
    10'b0000001101,
    10'b0001011001,
    10'b0100001101,
    10'b0010011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000011110,
    10'b0010000111,
    10'b0000000000,
    10'b0111000100,
    10'b0110001000,
    10'b1000010000,
    10'b0010000000,
    10'b0101011000,
    10'b0101100100,
    10'b0100011000,
    10'b1001100001,
    10'b0001000101,
    10'b0100100101,
    10'b1000011001,
    10'b0100001001,
    10'b0111001001,
    10'b1001011101,
    10'b0100100001,
    10'b0000010101,
    10'b0111011101,
    10'b0000001001,
    10'b0000011101,
    10'b0001100101,
    10'b0010001101,
    10'b0101010101,
    10'b0011011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0001001011,
    10'b1001011000,
    10'b0110001000,
    10'b0011100100,
    10'b0110001100,
    10'b1001100100,
    10'b0101100100,
    10'b1000000100,
    10'b0000011100,
    10'b0100001000,
    10'b0001010000,
    10'b0011000100,
    10'b0110100100,
    10'b1000010000,
    10'b0011010100,
    10'b1000010100,
    10'b0101010000,
    10'b1000100001,
    10'b0000000101,
    10'b0010011101,
    10'b0111011101,
    10'b0100100101,
    10'b0111010101,
    10'b0000100101,
    10'b0101001101,
    10'b0000010001,
    10'b1001010101,
    10'b0111001001,
    10'b0101000101,
    10'b1111111100,
    10'b1111111100,
    10'b0001001010,
    10'b0111100011,
    10'b0111100100,
    10'b0000100000,
    10'b0011100000,
    10'b0100100100,
    10'b1001001100,
    10'b0100000100,
    10'b0011011100,
    10'b1000000100,
    10'b0111010000,
    10'b0110011100,
    10'b0010011000,
    10'b1001011000,
    10'b0010000101,
    10'b1000100101,
    10'b0100100001,
    10'b0010010001,
    10'b0000000001,
    10'b0001011001,
    10'b0001001101,
    10'b0110100101,
    10'b1000100001,
    10'b0011001101,
    10'b0001000101,
    10'b0000011101,
    10'b0010100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111000110,
    10'b0001100011,
    10'b0101000000,
    10'b1000001100,
    10'b0100011100,
    10'b0111000000,
    10'b0111011100,
    10'b0001001100,
    10'b0101011100,
    10'b0011100000,
    10'b0110011100,
    10'b0011001000,
    10'b0100100100,
    10'b0110100000,
    10'b0001001000,
    10'b1000000101,
    10'b0010011101,
    10'b0100000001,
    10'b0000001001,
    10'b0010010001,
    10'b0000100101,
    10'b0011100101,
    10'b0101100001,
    10'b0011000001,
    10'b0100000101,
    10'b1001000001,
    10'b0100010101,
    10'b1001010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0001000111,
    10'b0100001100,
    10'b1001100000,
    10'b0101100100,
    10'b0001000000,
    10'b0001100100,
    10'b0100001000,
    10'b1001001000,
    10'b0111001000,
    10'b1001010100,
    10'b1000000000,
    10'b0110011100,
    10'b0100100100,
    10'b0101001000,
    10'b0110100101,
    10'b0010000101,
    10'b0011010001,
    10'b1000100101,
    10'b0010000001,
    10'b0011100001,
    10'b0011000101,
    10'b0001010101,
    10'b0000010101,
    10'b0001001001,
    10'b0100011001,
    10'b0001010001,
    10'b0101100001,
    10'b0101000001,
    10'b1001000001,
    10'b1000010101,
    10'b1000001001,
    10'b0001100010,
    10'b0111000111,
    10'b0000100100,
    10'b0100001100,
    10'b0001000100,
    10'b0010010100,
    10'b0011000000,
    10'b0000001100,
    10'b1000100000,
    10'b0101000000,
    10'b0001000000,
    10'b0011001000,
    10'b0000100001,
    10'b0110000001,
    10'b0110010101,
    10'b0110000101,
    10'b1001001101,
    10'b0001001101,
    10'b0101000101,
    10'b0100011001,
    10'b1001100001,
    10'b1001100101,
    10'b0111011001,
    10'b0000011101,
    10'b0101011001,
    10'b0111000001,
    10'b0100010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0011000110,
    10'b1000100011,
    10'b0000100000,
    10'b0011001100,
    10'b0011011100,
    10'b0011010000,
    10'b0110001100,
    10'b0010001000,
    10'b1001001100,
    10'b0000000000,
    10'b0010100100,
    10'b0000010000,
    10'b1001011000,
    10'b0011000000,
    10'b0100000101,
    10'b1000100101,
    10'b0010000001,
    10'b0010100001,
    10'b0100100101,
    10'b0100001001,
    10'b0000011101,
    10'b0001010001,
    10'b0111011101,
    10'b0100011101,
    10'b0010001101,
    10'b1000000001,
    10'b0101001101,
    10'b0101011001,
    10'b0100100001,
    10'b0100010101,
    10'b0010000101,
    10'b0111100001,
    10'b0010100010,
    10'b1000001011,
    10'b0000010100,
    10'b0111100100,
    10'b0110001000,
    10'b0101011000,
    10'b1001011100,
    10'b0100010000,
    10'b0101100100,
    10'b0111000000,
    10'b0110100100,
    10'b0010011100,
    10'b0110001100,
    10'b0001100001,
    10'b1001001001,
    10'b0101100001,
    10'b0010010101,
    10'b0011010101,
    10'b0010000001,
    10'b1001000101,
    10'b1001000001,
    10'b0101010001,
    10'b0100000101,
    10'b0100001101,
    10'b0001001101,
    10'b0001000001,
    10'b0011100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0101000100,
    10'b0110010000,
    10'b0000100100,
    10'b0110011100,
    10'b0111001000,
    10'b0111010000,
    10'b0101000000,
    10'b1000000000,
    10'b0111100100,
    10'b0101011000,
    10'b1001100001,
    10'b0000001101,
    10'b0111001101,
    10'b0000001001,
    10'b0110001101,
    10'b1000100101,
    10'b1000010101,
    10'b1001001101,
    10'b1001011001,
    10'b0001011101,
    10'b0000010001,
    10'b0010010101,
    10'b0011011001,
    10'b0001100101,
    10'b0011000101,
    10'b0110100101,
    10'b0011100101,
    10'b1001000001,
    10'b0010100101,
    10'b1111111100,
    10'b0001000110,
    10'b1000011111,
    10'b0011100000,
    10'b1001010100,
    10'b0000100000,
    10'b1001011100,
    10'b0001010000,
    10'b0001100100,
    10'b0100010000,
    10'b0010011000,
    10'b0111010100,
    10'b0110000100,
    10'b0100011000,
    10'b0100011100,
    10'b0100000100,
    10'b0011000000,
    10'b0001000001,
    10'b1001011101,
    10'b0100010101,
    10'b0100100001,
    10'b0001001001,
    10'b0000001101,
    10'b0011011101,
    10'b0010100101,
    10'b0110001001,
    10'b0000010001,
    10'b0010001001,
    10'b0101010001,
    10'b0101001101,
    10'b0001001101,
    10'b0110010101,
    10'b1111111100,
    10'b0110000110,
    10'b0001100011,
    10'b0001000100,
    10'b0100010100,
    10'b0000011100,
    10'b0000000000,
    10'b0011100000,
    10'b0001100100,
    10'b0010000100,
    10'b1000000000,
    10'b0111001000,
    10'b0111001001,
    10'b0001011101,
    10'b1001000101,
    10'b0111001101,
    10'b1001100101,
    10'b0001001101,
    10'b0010010101,
    10'b0000010101,
    10'b0110011001,
    10'b0011010001,
    10'b0010100101,
    10'b1001010001,
    10'b0011001001,
    10'b0101000001,
    10'b1000001001,
    10'b0110010001,
    10'b0100100001,
    10'b0111000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000011110,
    10'b0001001011,
    10'b0010000100,
    10'b0000100000,
    10'b0110011000,
    10'b0100011000,
    10'b0101010000,
    10'b0000010100,
    10'b0001100000,
    10'b1001000100,
    10'b1001100000,
    10'b0111100001,
    10'b0000001001,
    10'b0001010001,
    10'b1001010001,
    10'b0110001101,
    10'b0000000001,
    10'b0010010001,
    10'b0001001101,
    10'b0100001001,
    10'b1000001101,
    10'b0100000001,
    10'b0010000001,
    10'b0111010101,
    10'b0111001001,
    10'b0011001001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0001000111,
    10'b0111011100,
    10'b1001011100,
    10'b0101001000,
    10'b1001011000,
    10'b0100001100,
    10'b0010011100,
    10'b0110011100,
    10'b0101010000,
    10'b0111011000,
    10'b1001100100,
    10'b1001001000,
    10'b0111001100,
    10'b0011011000,
    10'b0011010000,
    10'b0000010000,
    10'b0110100001,
    10'b0000001001,
    10'b1000010101,
    10'b0010000101,
    10'b0111000001,
    10'b0011000001,
    10'b0110001001,
    10'b0000000001,
    10'b0000001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001110,
    10'b0001100011,
    10'b1000100000,
    10'b0100001100,
    10'b0111000100,
    10'b0100011100,
    10'b0011001100,
    10'b1001000000,
    10'b0110001000,
    10'b0110010000,
    10'b0101001000,
    10'b0111001101,
    10'b0000011101,
    10'b0110011101,
    10'b0110010101,
    10'b1001100101,
    10'b0000000101,
    10'b0101011001,
    10'b0111100001,
    10'b1000011101,
    10'b0000100001,
    10'b0101100001,
    10'b1000010001,
    10'b0111000001,
    10'b0100000101,
    10'b0111010101,
    10'b0001001101,
    10'b0101011101,
    10'b1001000101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0010011111,
    10'b0110100000,
    10'b0011010100,
    10'b1001011100,
    10'b0100010100,
    10'b0100010000,
    10'b0101000100,
    10'b1001011000,
    10'b1000011100,
    10'b0000010000,
    10'b0000010100,
    10'b0000100000,
    10'b0000000100,
    10'b0010000000,
    10'b0100000000,
    10'b0010100000,
    10'b0010010000,
    10'b1001000100,
    10'b0011000000,
    10'b1000001001,
    10'b0001011001,
    10'b0001010001,
    10'b0101011001,
    10'b0100000101,
    10'b0001100101,
    10'b0111010001,
    10'b0111100001,
    10'b0001010101,
    10'b1000011001,
    10'b1000001101,
    10'b1111111100,
    10'b1000100010,
    10'b0010000111,
    10'b0110100000,
    10'b0000100100,
    10'b1000000000,
    10'b0000010100,
    10'b1001001100,
    10'b0000010000,
    10'b0010011100,
    10'b0011100000,
    10'b0001001100,
    10'b1000010000,
    10'b0111100101,
    10'b0011000001,
    10'b0110001101,
    10'b0001010001,
    10'b0111011101,
    10'b0110011101,
    10'b0011010101,
    10'b0111000001,
    10'b0111001001,
    10'b0101001001,
    10'b0110100101,
    10'b0100100101,
    10'b0110000001,
    10'b0000011001,
    10'b0100100001,
    10'b0111010001,
    10'b0011001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000001011,
    10'b0011010100,
    10'b1001011100,
    10'b0100000000,
    10'b0001000100,
    10'b0100100000,
    10'b0110010000,
    10'b0011011000,
    10'b0011001100,
    10'b0111100100,
    10'b0010000100,
    10'b0000000100,
    10'b0011000100,
    10'b0001011101,
    10'b1000000101,
    10'b0000011001,
    10'b0011100101,
    10'b1000011101,
    10'b0000000001,
    10'b0110011101,
    10'b0010001101,
    10'b0001011001,
    10'b0001100101,
    10'b0110001101,
    10'b0110000001,
    10'b0100000101,
    10'b0101011101,
    10'b0010010001,
    10'b0000010101,
    10'b0000010001,
    10'b1111111100,
    10'b1000001010,
    10'b0010100011,
    10'b0110100100,
    10'b1000000100,
    10'b0110001000,
    10'b0010000000,
    10'b0010001100,
    10'b0010010100,
    10'b0110011100,
    10'b0101100100,
    10'b0111100000,
    10'b0001011000,
    10'b0011000000,
    10'b0100000000,
    10'b0110011000,
    10'b1001001001,
    10'b0011100101,
    10'b0100100101,
    10'b0011011101,
    10'b1000011101,
    10'b1000100001,
    10'b1000001101,
    10'b0011010101,
    10'b0100000101,
    10'b1001000101,
    10'b0111100101,
    10'b0110000101,
    10'b0111001001,
    10'b0000100001,
    10'b1000000001,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b1000011111,
    10'b0010100100,
    10'b0011001000,
    10'b0010001100,
    10'b1001000100,
    10'b0101000000,
    10'b1001001000,
    10'b1000010000,
    10'b0011000000,
    10'b0010000000,
    10'b0110001000,
    10'b1000001000,
    10'b0101011100,
    10'b0010000001,
    10'b1000011001,
    10'b1001010101,
    10'b0101011001,
    10'b0000011101,
    10'b0001001101,
    10'b0100010101,
    10'b0010011001,
    10'b0111000001,
    10'b0101010101,
    10'b1001100001,
    10'b0001100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001100011,
    10'b0101100100,
    10'b0100011000,
    10'b0000011000,
    10'b0101010100,
    10'b1001010100,
    10'b0010000000,
    10'b0111001100,
    10'b1000011000,
    10'b1001001000,
    10'b0111000000,
    10'b0110010000,
    10'b0111000100,
    10'b0111001001,
    10'b0000100001,
    10'b0001010001,
    10'b0010010101,
    10'b0011000001,
    10'b0111010001,
    10'b0011100001,
    10'b1001000101,
    10'b0011011001,
    10'b0110001001,
    10'b0101000001,
    10'b0110100101,
    10'b0000100101,
    10'b0101010001,
    10'b0000010101,
    10'b1000010001,
    10'b0111100001,
    10'b0110100001,
    10'b0011000110,
    10'b1000100011,
    10'b1000001000,
    10'b0010001100,
    10'b0001011100,
    10'b0010000000,
    10'b0100011100,
    10'b0100010100,
    10'b0011001100,
    10'b0000011000,
    10'b0110011100,
    10'b0000011100,
    10'b1000001100,
    10'b0010000001,
    10'b1001100001,
    10'b0111000001,
    10'b0011001001,
    10'b0000001101,
    10'b0011010001,
    10'b1001011101,
    10'b0110001001,
    10'b0101010001,
    10'b0100001001,
    10'b0110100001,
    10'b0001011001,
    10'b0010010101,
    10'b0001000101,
    10'b0010010001,
    10'b0011100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111001010,
    10'b0001100011,
    10'b0000001100,
    10'b1001001100,
    10'b1000100000,
    10'b0100001000,
    10'b0111011100,
    10'b0000100000,
    10'b0001001000,
    10'b0001100100,
    10'b0110001100,
    10'b0011001100,
    10'b1001001000,
    10'b0111000000,
    10'b0110011100,
    10'b1001011100,
    10'b0110100100,
    10'b0110000101,
    10'b0000100001,
    10'b0011000101,
    10'b1000001101,
    10'b0000010101,
    10'b0101010101,
    10'b0000011001,
    10'b0101011101,
    10'b0101001001,
    10'b0101010001,
    10'b0111100001,
    10'b1000001001,
    10'b1000010001,
    10'b0001011001,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0001000000,
    10'b0110100100,
    10'b0011000000,
    10'b0101011000,
    10'b0101001000,
    10'b1000011000,
    10'b1000000100,
    10'b1001010000,
    10'b0101100000,
    10'b1001000100,
    10'b1001100000,
    10'b0111011100,
    10'b0011100000,
    10'b0101000000,
    10'b0100011000,
    10'b0100011100,
    10'b1001100101,
    10'b0000001101,
    10'b0011000101,
    10'b0110010001,
    10'b0010001001,
    10'b0100010101,
    10'b1001011101,
    10'b0100001001,
    10'b0000000101,
    10'b1001000001,
    10'b0110011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001011110,
    10'b1000001011,
    10'b0000000100,
    10'b0001000000,
    10'b0101010100,
    10'b0010001100,
    10'b0100000000,
    10'b0010100100,
    10'b0100000100,
    10'b1001100100,
    10'b0110011100,
    10'b0111010100,
    10'b0100100100,
    10'b1000010000,
    10'b1000011100,
    10'b0010000000,
    10'b0001010000,
    10'b0111000000,
    10'b0101000000,
    10'b0100001000,
    10'b0000011101,
    10'b1000001101,
    10'b0111001001,
    10'b0101100101,
    10'b1000100001,
    10'b0001001001,
    10'b0010011101,
    10'b1000100101,
    10'b1001000001,
    10'b1001010101,
    10'b0101100001,
    10'b0101001001,
    10'b0111100010,
    10'b0001000111,
    10'b0011011100,
    10'b0100001100,
    10'b0011001000,
    10'b0001010000,
    10'b0001001100,
    10'b1000011000,
    10'b0011001100,
    10'b1001000000,
    10'b0111100100,
    10'b0001010100,
    10'b0101011100,
    10'b0001011100,
    10'b1001011100,
    10'b1000100000,
    10'b0000000000,
    10'b0001000000,
    10'b0111011101,
    10'b0000001001,
    10'b0010011001,
    10'b0010010101,
    10'b0111000001,
    10'b0001001001,
    10'b0010000001,
    10'b1001100001,
    10'b0110011101,
    10'b0100011001,
    10'b0000000101,
    10'b0101010101,
    10'b1111111100,
    10'b1111111100,
    10'b0111011110,
    10'b0001000111,
    10'b0001001100,
    10'b0010100000,
    10'b0000010000,
    10'b0100001100,
    10'b1000011000,
    10'b1000001100,
    10'b0100010000,
    10'b1001000100,
    10'b0010000000,
    10'b0111010000,
    10'b0101011100,
    10'b0101000100,
    10'b0110001100,
    10'b0101100100,
    10'b0111000100,
    10'b1000011101,
    10'b0010000001,
    10'b0001001001,
    10'b0110100001,
    10'b1001010001,
    10'b0101001001,
    10'b0001000001,
    10'b1000001001,
    10'b0001011101,
    10'b1000000101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b0110100011,
    10'b0011000100,
    10'b0010000000,
    10'b0110000000,
    10'b0010010100,
    10'b0010011100,
    10'b0110100100,
    10'b0001001000,
    10'b0100001000,
    10'b0101100000,
    10'b0001001001,
    10'b0111100101,
    10'b0000001101,
    10'b0101010101,
    10'b0010100001,
    10'b0011100001,
    10'b1000001101,
    10'b0111000001,
    10'b0010100101,
    10'b1000000001,
    10'b1001010001,
    10'b0000000001,
    10'b0011001001,
    10'b0000000101,
    10'b0000100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111000110,
    10'b0001011111,
    10'b0111011100,
    10'b0011100100,
    10'b0101100100,
    10'b0101100000,
    10'b0111100000,
    10'b1000010100,
    10'b0100100000,
    10'b0000100000,
    10'b0101001100,
    10'b1001001000,
    10'b0001010000,
    10'b0000001100,
    10'b0011001100,
    10'b0001000000,
    10'b0011000000,
    10'b0111001001,
    10'b0010011001,
    10'b0100010001,
    10'b0101010101,
    10'b0011010101,
    10'b0100001001,
    10'b0101000001,
    10'b0111001101,
    10'b0010010101,
    10'b0110100101,
    10'b1001100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111000110,
    10'b0001100011,
    10'b1000000100,
    10'b0010000000,
    10'b1000001100,
    10'b0101100100,
    10'b0001000000,
    10'b0001001000,
    10'b0100001000,
    10'b0110010000,
    10'b0111100100,
    10'b0100100000,
    10'b1000000000,
    10'b0010100000,
    10'b1001000000,
    10'b0110000001,
    10'b0010011101,
    10'b0110000101,
    10'b0000100001,
    10'b1001011101,
    10'b0011100101,
    10'b1001100101,
    10'b0100100101,
    10'b1000011001,
    10'b0100010001,
    10'b0100010101,
    10'b0100011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b1000100011,
    10'b1000011000,
    10'b1000011100,
    10'b0010000000,
    10'b0010001000,
    10'b0110010100,
    10'b1000010000,
    10'b1001011000,
    10'b0100011000,
    10'b0111100100,
    10'b0111011100,
    10'b0101001000,
    10'b1001011100,
    10'b0111000000,
    10'b0000100000,
    10'b0011100100,
    10'b0101001100,
    10'b0010001001,
    10'b1001100101,
    10'b0001100101,
    10'b0010011001,
    10'b0000011001,
    10'b0111010001,
    10'b0001011001,
    10'b0111000101,
    10'b0010001101,
    10'b0000010101,
    10'b0101100101,
    10'b0001100001,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0011100011,
    10'b0101001100,
    10'b0001000100,
    10'b0110100000,
    10'b1000011100,
    10'b0100001000,
    10'b1000100000,
    10'b0110011100,
    10'b0111100100,
    10'b0111000100,
    10'b0111001000,
    10'b0101001000,
    10'b0000011000,
    10'b0111000001,
    10'b0011011101,
    10'b0100000101,
    10'b0010000001,
    10'b0001100101,
    10'b0000010001,
    10'b1001010101,
    10'b0011011001,
    10'b0110001101,
    10'b0001010001,
    10'b1001001101,
    10'b0001000001,
    10'b0001001101,
    10'b0111010001,
    10'b0010001001,
    10'b1001000101,
    10'b1111111100,
    10'b1111111100,
    10'b0001011110,
    10'b1000000111,
    10'b1001001000,
    10'b0101100100,
    10'b0101011100,
    10'b0100001000,
    10'b0110000100,
    10'b1000000000,
    10'b0100100000,
    10'b1000100000,
    10'b1001001100,
    10'b0000011101,
    10'b0111001001,
    10'b0100011001,
    10'b1000001101,
    10'b0110010001,
    10'b0111010001,
    10'b1001100101,
    10'b0100001101,
    10'b0000010101,
    10'b0110000001,
    10'b0111100101,
    10'b0000000001,
    10'b0100100101,
    10'b0011010101,
    10'b0010011101,
    10'b0110010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000001111,
    10'b0011001100,
    10'b0010010000,
    10'b0001010000,
    10'b0000001000,
    10'b1000011000,
    10'b0110000100,
    10'b0010011000,
    10'b0000100000,
    10'b1001011000,
    10'b0011010000,
    10'b0010000000,
    10'b0111011100,
    10'b1001010100,
    10'b0111100100,
    10'b0011010100,
    10'b1001001000,
    10'b0001000000,
    10'b0000000000,
    10'b1001011100,
    10'b0000011101,
    10'b1001001101,
    10'b0011100001,
    10'b0110010001,
    10'b0000010101,
    10'b1001100001,
    10'b0111010101,
    10'b0111010001,
    10'b0110011001,
    10'b0111000101,
    10'b1001000101,
    10'b0001000110,
    10'b1000011011,
    10'b0001100000,
    10'b0000001100,
    10'b0010100100,
    10'b1001010100,
    10'b0010000000,
    10'b0101100100,
    10'b0111010000,
    10'b0101001000,
    10'b0101001100,
    10'b0000000000,
    10'b0000100000,
    10'b0110100000,
    10'b0111000100,
    10'b0001000000,
    10'b0000000001,
    10'b1001011001,
    10'b0101100001,
    10'b0010001101,
    10'b0000011001,
    10'b0100100101,
    10'b0001010101,
    10'b0011000001,
    10'b1001001001,
    10'b0000011101,
    10'b0101010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001110,
    10'b0001100011,
    10'b0001000000,
    10'b0111100100,
    10'b1001100100,
    10'b0010010000,
    10'b1000100100,
    10'b0101010000,
    10'b0101100000,
    10'b0110100100,
    10'b0010001000,
    10'b1001010001,
    10'b0001100101,
    10'b0000010101,
    10'b0100001001,
    10'b0101001001,
    10'b1000011001,
    10'b0111001001,
    10'b0010100101,
    10'b0011011001,
    10'b0111000001,
    10'b0101011101,
    10'b0100000001,
    10'b0000100001,
    10'b0000011001,
    10'b1000010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0001000111,
    10'b1001001100,
    10'b0111011000,
    10'b1000100000,
    10'b0100001100,
    10'b0010000100,
    10'b0110100000,
    10'b0101100100,
    10'b0101000000,
    10'b0110000000,
    10'b0011010100,
    10'b0100000100,
    10'b0110001000,
    10'b0100000000,
    10'b0011100000,
    10'b0110011101,
    10'b0010000001,
    10'b0010001101,
    10'b0000011001,
    10'b0100011101,
    10'b0010011001,
    10'b1001000001,
    10'b0100010001,
    10'b1001011001,
    10'b0001010001,
    10'b0111100101,
    10'b0011100101,
    10'b0011001001,
    10'b1000001001,
    10'b0011010001,
    10'b0111010101,
    10'b0110100010,
    10'b0001000111,
    10'b0110011100,
    10'b0101010000,
    10'b0000100100,
    10'b1000000000,
    10'b1001001000,
    10'b1000000100,
    10'b0010011100,
    10'b0100000000,
    10'b0001011100,
    10'b0101001100,
    10'b0010010000,
    10'b1000011100,
    10'b1001011100,
    10'b0111011101,
    10'b0000001001,
    10'b0011011001,
    10'b0101000101,
    10'b1001010001,
    10'b0111100101,
    10'b0010001101,
    10'b0011010101,
    10'b0011100101,
    10'b0011001001,
    10'b0001010001,
    10'b0011010001,
    10'b0001001101,
    10'b0000011001,
    10'b0001100001,
    10'b1000010101,
    10'b0010100001,
    10'b1000000110,
    10'b0011100011,
    10'b0000001000,
    10'b1001100000,
    10'b0000011100,
    10'b0111011100,
    10'b0000010000,
    10'b0000000100,
    10'b1000001100,
    10'b0101100000,
    10'b1001100100,
    10'b0001011100,
    10'b0001010000,
    10'b0001001100,
    10'b0111000101,
    10'b0010100001,
    10'b0011001101,
    10'b1001010001,
    10'b1000011101,
    10'b0011011001,
    10'b0111011001,
    10'b0001100101,
    10'b1001001101,
    10'b0011010101,
    10'b0111000001,
    10'b0010010101,
    10'b1001001001,
    10'b0100001001,
    10'b0111010101,
    10'b1001000101,
    10'b0100001101,
    10'b0101000101,
    10'b0010100010,
    10'b1000001011,
    10'b0101011100,
    10'b0000000100,
    10'b0000001000,
    10'b1001010100,
    10'b1000100100,
    10'b0001000100,
    10'b0010011100,
    10'b0110100000,
    10'b0000100000,
    10'b0011100100,
    10'b0110011100,
    10'b0101001000,
    10'b0111011100,
    10'b0100001100,
    10'b0011001000,
    10'b0011010000,
    10'b1001010000,
    10'b0010100101,
    10'b0111001101,
    10'b0011010101,
    10'b0000010001,
    10'b0100011101,
    10'b1000000001,
    10'b1000010101,
    10'b0010010101,
    10'b1001100101,
    10'b0011001101,
    10'b0010011001,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0000010100,
    10'b0100100100,
    10'b1000001100,
    10'b0010100000,
    10'b0011100000,
    10'b0101001000,
    10'b0011001000,
    10'b0110001100,
    10'b0110001000,
    10'b0101011000,
    10'b1001001100,
    10'b0110100000,
    10'b0001000100,
    10'b0111011101,
    10'b0010010001,
    10'b0000011101,
    10'b1000011001,
    10'b0010011101,
    10'b0110010101,
    10'b0100001101,
    10'b1001010101,
    10'b1001100001,
    10'b0111000001,
    10'b0001011101,
    10'b1001011101,
    10'b0011001101,
    10'b0111010001,
    10'b0100011101,
    10'b1000011101,
    10'b1111111100,
    10'b0001011110,
    10'b1000000111,
    10'b0010000000,
    10'b0110010000,
    10'b0000011100,
    10'b0101011000,
    10'b0011100100,
    10'b1000000000,
    10'b0010011100,
    10'b0011010100,
    10'b0011000100,
    10'b0001100100,
    10'b0011011100,
    10'b0110100000,
    10'b0000011001,
    10'b0111001001,
    10'b1001001101,
    10'b0110000001,
    10'b1001010101,
    10'b1000011001,
    10'b0000100001,
    10'b0100010101,
    10'b0011011001,
    10'b0011010001,
    10'b0100010001,
    10'b1001011001,
    10'b0001010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b0111001011,
    10'b1000100000,
    10'b0110011100,
    10'b0010001000,
    10'b0001001000,
    10'b0101100100,
    10'b0101010000,
    10'b0101001000,
    10'b0111100000,
    10'b0000001000,
    10'b0111011100,
    10'b1001011000,
    10'b1000001000,
    10'b0010011000,
    10'b0011000000,
    10'b0001100101,
    10'b0111001101,
    10'b0100000001,
    10'b0101100001,
    10'b0100001001,
    10'b0100100001,
    10'b0011100001,
    10'b0010000001,
    10'b0110001101,
    10'b0011001001,
    10'b0111000101,
    10'b1000011101,
    10'b0100010101,
    10'b1000011001,
    10'b0001001101,
    10'b1111111100,
    10'b0011000110,
    10'b1000100011,
    10'b0111000000,
    10'b0100100100,
    10'b0100000100,
    10'b0111011000,
    10'b1001000000,
    10'b0100001100,
    10'b0010000000,
    10'b1001010100,
    10'b0110000000,
    10'b1001100000,
    10'b0010010100,
    10'b0001001000,
    10'b0111000100,
    10'b0000000000,
    10'b0001011100,
    10'b1001011000,
    10'b0101001000,
    10'b0010001100,
    10'b0010000100,
    10'b0010000001,
    10'b0111100101,
    10'b1000011001,
    10'b0000001001,
    10'b0010011001,
    10'b0010011101,
    10'b0000000101,
    10'b0001000101,
    10'b0000100101,
    10'b0100010001,
    10'b0001000001,
    10'b1000000110,
    10'b0001100011,
    10'b0000000000,
    10'b0100100100,
    10'b1001011100,
    10'b0010010000,
    10'b0000011000,
    10'b1000100000,
    10'b0110011000,
    10'b0001001100,
    10'b0001000100,
    10'b0010000100,
    10'b0011001000,
    10'b1001100100,
    10'b0101001100,
    10'b1001010100,
    10'b1000100100,
    10'b0011100000,
    10'b0101000100,
    10'b0011010100,
    10'b1001000101,
    10'b0010011101,
    10'b0111001001,
    10'b0101011101,
    10'b0111010101,
    10'b0010001101,
    10'b1000011001,
    10'b0110100101,
    10'b0101100001,
    10'b0011000101,
    10'b0100010001,
    10'b0110010001,
    10'b1000100010,
    10'b0001001111,
    10'b0010011100,
    10'b0111001000,
    10'b0010010100,
    10'b0101000100,
    10'b0010010000,
    10'b0110011100,
    10'b0110100100,
    10'b0000100100,
    10'b0111011101,
    10'b0000010001,
    10'b1000011101,
    10'b0000000101,
    10'b1000000001,
    10'b0001010101,
    10'b1001011001,
    10'b0011001101,
    10'b0010011001,
    10'b0010100001,
    10'b0111100001,
    10'b0111010001,
    10'b0110100001,
    10'b0101000001,
    10'b0000011101,
    10'b0000010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b0111001011,
    10'b0111000100,
    10'b0100100100,
    10'b0000001100,
    10'b0110011100,
    10'b0000010100,
    10'b0111011100,
    10'b1000011100,
    10'b1001000000,
    10'b0010001000,
    10'b0010000100,
    10'b0111011000,
    10'b1001010100,
    10'b0001010000,
    10'b0100000000,
    10'b0010100101,
    10'b0111001101,
    10'b0100011101,
    10'b0110010001,
    10'b0000000101,
    10'b1001011101,
    10'b1001010001,
    10'b1000010001,
    10'b1000010101,
    10'b0111100001,
    10'b0010011101,
    10'b0000001001,
    10'b0111100101,
    10'b1000100101,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000100011,
    10'b0001010000,
    10'b0101000000,
    10'b0101010100,
    10'b0110010100,
    10'b1000000100,
    10'b1000011000,
    10'b0101001100,
    10'b1001100100,
    10'b0011011100,
    10'b0100000000,
    10'b0111100100,
    10'b0011000000,
    10'b0001000001,
    10'b0111100001,
    10'b0111011101,
    10'b0011011001,
    10'b0011001101,
    10'b0110100001,
    10'b1001010101,
    10'b1000001101,
    10'b0000011001,
    10'b0010001101,
    10'b0110011001,
    10'b1001001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001001110,
    10'b1000100011,
    10'b0101000100,
    10'b0100100000,
    10'b0110000100,
    10'b0001010100,
    10'b0100100100,
    10'b0100001100,
    10'b0001001000,
    10'b0010011000,
    10'b0101000000,
    10'b0010001000,
    10'b0001100000,
    10'b0100000100,
    10'b0110010100,
    10'b1001000100,
    10'b0110011000,
    10'b0001010001,
    10'b1000100101,
    10'b0111010001,
    10'b1000000101,
    10'b0111010101,
    10'b1001001101,
    10'b0010010101,
    10'b0001000101,
    10'b1000001001,
    10'b0110100101,
    10'b0111011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0110000110,
    10'b0001100011,
    10'b1000010100,
    10'b0101100100,
    10'b0011000000,
    10'b0010000100,
    10'b0000011000,
    10'b1001001000,
    10'b0111010100,
    10'b1000100000,
    10'b0011100100,
    10'b0000000000,
    10'b1001100100,
    10'b0111000000,
    10'b0100100000,
    10'b0111001001,
    10'b0000011101,
    10'b0110001001,
    10'b0101010101,
    10'b0000001101,
    10'b0010001101,
    10'b1000011001,
    10'b0110011001,
    10'b0100011001,
    10'b0001011001,
    10'b0001001101,
    10'b0011001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0010000111,
    10'b0111001100,
    10'b1000000100,
    10'b1000011000,
    10'b0010100100,
    10'b1000100000,
    10'b0100011000,
    10'b0001010000,
    10'b0111001000,
    10'b0100011100,
    10'b0010001100,
    10'b1001010000,
    10'b1001000000,
    10'b0111000000,
    10'b0001000000,
    10'b0110001000,
    10'b0110100100,
    10'b1000100101,
    10'b0001000001,
    10'b0000001001,
    10'b0000010001,
    10'b0010100001,
    10'b0001011001,
    10'b0110010101,
    10'b0000000101,
    10'b0000100001,
    10'b0001100001,
    10'b0101001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000100011,
    10'b0110011000,
    10'b0101011100,
    10'b1000011100,
    10'b1000000100,
    10'b1000001000,
    10'b0010001100,
    10'b0101010100,
    10'b1001100000,
    10'b0001000000,
    10'b0110000000,
    10'b0101001000,
    10'b1000001100,
    10'b1000100100,
    10'b0011000101,
    10'b0111100101,
    10'b0101010001,
    10'b0001100001,
    10'b0110010001,
    10'b0111011101,
    10'b0010010101,
    10'b0100010101,
    10'b0010011001,
    10'b0110011101,
    10'b0001010101,
    10'b0011000001,
    10'b0010100101,
    10'b0011010101,
    10'b0010001001,
    10'b0101000101,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0110001100,
    10'b0100011100,
    10'b0110100100,
    10'b0101100000,
    10'b0010100000,
    10'b0101010000,
    10'b0111001000,
    10'b0100001000,
    10'b0110100000,
    10'b0001000100,
    10'b0000010000,
    10'b0100000000,
    10'b0010001100,
    10'b0110011100,
    10'b0111011101,
    10'b0010001001,
    10'b1001100001,
    10'b0100000101,
    10'b0010011001,
    10'b0111100001,
    10'b0011010001,
    10'b0011011101,
    10'b0011000101,
    10'b0001100101,
    10'b1001000101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0010000111,
    10'b0011011100,
    10'b0000000000,
    10'b0011011000,
    10'b0001100000,
    10'b0100011100,
    10'b0001100100,
    10'b0011010000,
    10'b1001011100,
    10'b0001000000,
    10'b0001010100,
    10'b0000000100,
    10'b1001010000,
    10'b0010010100,
    10'b0000010000,
    10'b0100100100,
    10'b0011000000,
    10'b1000100001,
    10'b0011000101,
    10'b1000000001,
    10'b0100001001,
    10'b0100000001,
    10'b0011100101,
    10'b0011010101,
    10'b0001001001,
    10'b1000010101,
    10'b0000010101,
    10'b0001001101,
    10'b0111011001,
    10'b1111111100,
    10'b1111111100,
    10'b0110000110,
    10'b0001100011,
    10'b0110011100,
    10'b0100011000,
    10'b0010100100,
    10'b0010011100,
    10'b0111001000,
    10'b0101011000,
    10'b0110001100,
    10'b0101100100,
    10'b0010010100,
    10'b0110100000,
    10'b0001000000,
    10'b0100010100,
    10'b0101001001,
    10'b0000100001,
    10'b0010010001,
    10'b0011011101,
    10'b0011011001,
    10'b1001011101,
    10'b1000011001,
    10'b0011010001,
    10'b0011001101,
    10'b1001001101,
    10'b1000100101,
    10'b0110001001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001100011,
    10'b1001100100,
    10'b0010100100,
    10'b0001001100,
    10'b0101001100,
    10'b0001100100,
    10'b0011100000,
    10'b0010010000,
    10'b0101010100,
    10'b0111010000,
    10'b1000100000,
    10'b0000011000,
    10'b0011100100,
    10'b1001000101,
    10'b0001011101,
    10'b1001010101,
    10'b0110011101,
    10'b0100011001,
    10'b0001011001,
    10'b0110000001,
    10'b0011011101,
    10'b0111100101,
    10'b0101001001,
    10'b1001000001,
    10'b0110001001,
    10'b1000011101,
    10'b0010011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001011111,
    10'b0011100000,
    10'b0000010100,
    10'b1000010100,
    10'b1000100100,
    10'b0111000100,
    10'b0100100000,
    10'b0100000000,
    10'b0010001000,
    10'b0000010000,
    10'b1001010100,
    10'b0111000101,
    10'b0010011001,
    10'b0101001001,
    10'b0011100101,
    10'b1000011101,
    10'b0010011101,
    10'b0010000001,
    10'b0001010101,
    10'b1001100001,
    10'b0010001101,
    10'b0100100101,
    10'b1000001001,
    10'b0011011001,
    10'b1000010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000011010,
    10'b0001000111,
    10'b0101000100,
    10'b0010011000,
    10'b0000100100,
    10'b0000010100,
    10'b0000010000,
    10'b0000000100,
    10'b0110011100,
    10'b0111011100,
    10'b1000010000,
    10'b1001011100,
    10'b1001010101,
    10'b0001001001,
    10'b0110011001,
    10'b1000001001,
    10'b0100001001,
    10'b0001010101,
    10'b0100011001,
    10'b1001001001,
    10'b0100000001,
    10'b0000001001,
    10'b0111010001,
    10'b0100100001,
    10'b1001000001,
    10'b0011010001,
    10'b0010010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0010100011,
    10'b0110001000,
    10'b1001100000,
    10'b0011010000,
    10'b0000000100,
    10'b1001000000,
    10'b0000011100,
    10'b0100010100,
    10'b0011000100,
    10'b1000011000,
    10'b0001011100,
    10'b0010010000,
    10'b0100000000,
    10'b0010011100,
    10'b0101100100,
    10'b0100011100,
    10'b1001000101,
    10'b0001100001,
    10'b0000010001,
    10'b1000011101,
    10'b0111010001,
    10'b0000100101,
    10'b0100000101,
    10'b0110000001,
    10'b0111100001,
    10'b0110100101,
    10'b0110011101,
    10'b0000100001,
    10'b1001010001,
    10'b1111111100,
    10'b1111111100,
    10'b0111001010,
    10'b0001100011,
    10'b0000000100,
    10'b0101000000,
    10'b0100000100,
    10'b1000001100,
    10'b1000010100,
    10'b0111100000,
    10'b0001001100,
    10'b1001001000,
    10'b0000001100,
    10'b0011100100,
    10'b1000010000,
    10'b0010001100,
    10'b0010000100,
    10'b1000001101,
    10'b0000011101,
    10'b1001000001,
    10'b0011010001,
    10'b0001000001,
    10'b1001010001,
    10'b0111000101,
    10'b0001000101,
    10'b0100010101,
    10'b0000100101,
    10'b0001010001,
    10'b0001010101,
    10'b0010000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0001000111,
    10'b0001100000,
    10'b0011100000,
    10'b0011010100,
    10'b0011011000,
    10'b0111001100,
    10'b0010010100,
    10'b1001001000,
    10'b0100010100,
    10'b0000010000,
    10'b0101100100,
    10'b1000010100,
    10'b0001010100,
    10'b1000100101,
    10'b0010000001,
    10'b0010001101,
    10'b0000100001,
    10'b0100100101,
    10'b0110001101,
    10'b0111000001,
    10'b0000011001,
    10'b0000001001,
    10'b1001011101,
    10'b0010011101,
    10'b0110011001,
    10'b0101000101,
    10'b0101011101,
    10'b0111011001,
    10'b0010100101,
    10'b1111111100,
    10'b1111111100,
    10'b0111001010,
    10'b0001100011,
    10'b0001000000,
    10'b0100000000,
    10'b0011011100,
    10'b0001011100,
    10'b0000010100,
    10'b0011001100,
    10'b0000000100,
    10'b0000011000,
    10'b0110100100,
    10'b1001001000,
    10'b0101011100,
    10'b0000011100,
    10'b1000000101,
    10'b0001011101,
    10'b0101001101,
    10'b0111001101,
    10'b0001000101,
    10'b0010001101,
    10'b0000010001,
    10'b0000100001,
    10'b0101100101,
    10'b0100100001,
    10'b1001100001,
    10'b0100001001,
    10'b0010000001,
    10'b0001001001,
    10'b0011010101,
    10'b0111100101,
    10'b0101011001,
    10'b1111111100,
    10'b0001011010,
    10'b1000000111,
    10'b0001000100,
    10'b0100010100,
    10'b0001001000,
    10'b0010000000,
    10'b0000100100,
    10'b0000011100,
    10'b0110010000,
    10'b0010011100,
    10'b0101010000,
    10'b1000000000,
    10'b1001011100,
    10'b1001000100,
    10'b0111011000,
    10'b0000010000,
    10'b0110011000,
    10'b0001010101,
    10'b0111000101,
    10'b0000000101,
    10'b0101100101,
    10'b0111001001,
    10'b0111001101,
    10'b0010100001,
    10'b1000001101,
    10'b1001001101,
    10'b0010000101,
    10'b0001100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010011110,
    10'b1000000111,
    10'b0101001000,
    10'b0010100100,
    10'b1001100000,
    10'b0001000000,
    10'b1000100000,
    10'b0111010000,
    10'b0110001000,
    10'b0001001100,
    10'b0000100000,
    10'b1000001000,
    10'b0000011000,
    10'b0001011101,
    10'b1001000001,
    10'b0000100101,
    10'b0110011001,
    10'b0111010101,
    10'b0010000101,
    10'b0010100001,
    10'b0111100101,
    10'b0001011001,
    10'b0010000001,
    10'b0100100101,
    10'b0110100101,
    10'b0111011101,
    10'b1001100101,
    10'b1001011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001001010,
    10'b1000100011,
    10'b1000100100,
    10'b1000001000,
    10'b1001011000,
    10'b0100010100,
    10'b0000100100,
    10'b1001000000,
    10'b0001001100,
    10'b0000001000,
    10'b0011000000,
    10'b0001011100,
    10'b0110000100,
    10'b0100100100,
    10'b0101001000,
    10'b0100010000,
    10'b0001001101,
    10'b1001100101,
    10'b0101011001,
    10'b0100000101,
    10'b0000100001,
    10'b0110000001,
    10'b1001001001,
    10'b0010000001,
    10'b0111001101,
    10'b0111100001,
    10'b0110100101,
    10'b0011001101,
    10'b1000010101,
    10'b0000011101,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000011111,
    10'b1001010100,
    10'b0000011100,
    10'b0101100000,
    10'b0010001100,
    10'b0010100100,
    10'b1000100000,
    10'b0110100100,
    10'b0011011100,
    10'b1001100000,
    10'b0001000000,
    10'b0110000100,
    10'b1000000100,
    10'b0001000001,
    10'b1000100001,
    10'b0000000001,
    10'b0000011001,
    10'b0011100001,
    10'b0100010001,
    10'b0000100101,
    10'b0011011001,
    10'b0010001001,
    10'b0000010001,
    10'b0001010001,
    10'b0100011001,
    10'b0110001001,
    10'b0001011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001011,
    10'b0010000100,
    10'b1001000100,
    10'b0110100000,
    10'b0110011000,
    10'b0100000100,
    10'b0101000000,
    10'b1000001000,
    10'b0110011100,
    10'b0000010000,
    10'b0110001100,
    10'b0001010100,
    10'b1000011000,
    10'b0001100000,
    10'b1001011100,
    10'b0111001100,
    10'b1001000000,
    10'b1001100001,
    10'b0010000101,
    10'b0101011001,
    10'b1000100101,
    10'b1001001101,
    10'b0000001101,
    10'b0001011001,
    10'b0111010101,
    10'b0000100001,
    10'b0011001101,
    10'b0100010001,
    10'b0111100001,
    10'b1000010101,
    10'b1001010101,
    10'b0010011110,
    10'b1000000111,
    10'b0110100000,
    10'b0000100000,
    10'b0100001100,
    10'b1000011100,
    10'b0010001000,
    10'b0111011000,
    10'b1001000000,
    10'b0001010000,
    10'b0000011100,
    10'b1001100000,
    10'b1001010100,
    10'b0011000000,
    10'b0101001000,
    10'b0001011001,
    10'b0111000001,
    10'b0011010101,
    10'b0011100001,
    10'b0001001101,
    10'b1001100101,
    10'b0000010001,
    10'b1001011001,
    10'b0010010101,
    10'b0101011001,
    10'b0110011101,
    10'b1000000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010001010,
    10'b1000100011,
    10'b0011100100,
    10'b1000001100,
    10'b0110001100,
    10'b1000010100,
    10'b0010000000,
    10'b0101001100,
    10'b1001000000,
    10'b0001000100,
    10'b1001010100,
    10'b0000100000,
    10'b0011100000,
    10'b0100100000,
    10'b0100001000,
    10'b0001001101,
    10'b1001100101,
    10'b0010100001,
    10'b0110011101,
    10'b0001010101,
    10'b0001100101,
    10'b0010001101,
    10'b1001000101,
    10'b0100011101,
    10'b0101010001,
    10'b0110010001,
    10'b0101100101,
    10'b0100000101,
    10'b0101011001,
    10'b0001010001,
    10'b1111111100,
    10'b1111111100,
    10'b0011100010,
    10'b1000000111,
    10'b0000010100,
    10'b0010000100,
    10'b0010100000,
    10'b1001001100,
    10'b1001000000,
    10'b0010011000,
    10'b0001000100,
    10'b0000010000,
    10'b1001000100,
    10'b0000001100,
    10'b0011001100,
    10'b0001100000,
    10'b0100011101,
    10'b1000000001,
    10'b0001011001,
    10'b1000011001,
    10'b0000001001,
    10'b0011010101,
    10'b0110001101,
    10'b0011000101,
    10'b0101100101,
    10'b1000001101,
    10'b1001100001,
    10'b0111011101,
    10'b0100100101,
    10'b0111000101,
    10'b0010011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b0111000111,
    10'b0011010000,
    10'b0010100100,
    10'b0001100100,
    10'b0111100100,
    10'b0000001100,
    10'b1000000000,
    10'b1001000000,
    10'b1001100100,
    10'b0101001100,
    10'b0110011000,
    10'b0011010100,
    10'b0000011101,
    10'b1000000101,
    10'b0101011001,
    10'b1000100101,
    10'b1001001101,
    10'b0001001101,
    10'b1000011101,
    10'b0110010001,
    10'b0101000101,
    10'b0100010101,
    10'b0110001001,
    10'b0010011101,
    10'b1001011101,
    10'b0001011101,
    10'b0000100101,
    10'b1000001101,
    10'b0010000101,
    10'b0010000001,
    10'b0001000001,
    10'b0001100010,
    10'b1000000111,
    10'b0110011100,
    10'b0111001100,
    10'b1000100000,
    10'b0000001100,
    10'b0101100100,
    10'b0111010100,
    10'b0011001000,
    10'b0000010000,
    10'b0101011100,
    10'b1001010000,
    10'b0010000000,
    10'b0101010100,
    10'b0100100000,
    10'b0110011000,
    10'b1001010100,
    10'b0001000100,
    10'b0001100101,
    10'b0111001001,
    10'b1001011101,
    10'b1001100101,
    10'b0011011001,
    10'b0101100001,
    10'b0001010101,
    10'b1001000001,
    10'b0111011001,
    10'b0100100101,
    10'b0011000001,
    10'b0110100101,
    10'b1111111100,
    10'b1111111100,
    10'b0111100010,
    10'b0010000111,
    10'b0110100100,
    10'b0001010000,
    10'b0000010100,
    10'b0001010100,
    10'b0110001100,
    10'b0100001000,
    10'b0000100000,
    10'b0000001000,
    10'b1000100000,
    10'b0100100100,
    10'b0000001100,
    10'b0101000000,
    10'b0100011100,
    10'b0011001000,
    10'b0000011000,
    10'b0001000100,
    10'b0110100001,
    10'b0001000001,
    10'b0010001101,
    10'b0100010001,
    10'b0001001101,
    10'b0010000001,
    10'b1001100001,
    10'b1001000001,
    10'b0101011101,
    10'b0111000101,
    10'b1001000101,
    10'b0101001101,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000100011,
    10'b0110011100,
    10'b0101100100,
    10'b0011000000,
    10'b0000001100,
    10'b0000011100,
    10'b0001100000,
    10'b0111100000,
    10'b0100001100,
    10'b0101011100,
    10'b0001011100,
    10'b1001010000,
    10'b0011001001,
    10'b1001100101,
    10'b0011100101,
    10'b0011010101,
    10'b0100000001,
    10'b0011001101,
    10'b0000000101,
    10'b0110100101,
    10'b0100000101,
    10'b0000001001,
    10'b1001000001,
    10'b1000010101,
    10'b1001000101,
    10'b0110011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b1000100011,
    10'b0011000100,
    10'b0001010100,
    10'b1001000100,
    10'b1000010100,
    10'b0010011000,
    10'b0111001000,
    10'b0000010100,
    10'b0001011000,
    10'b0111100100,
    10'b0110000100,
    10'b0110010000,
    10'b1000000000,
    10'b1001010100,
    10'b0111011000,
    10'b0101001100,
    10'b0110011000,
    10'b0000011100,
    10'b0001000001,
    10'b1000100101,
    10'b0001001001,
    10'b0000100101,
    10'b0110010101,
    10'b0101100101,
    10'b0011100001,
    10'b0010000001,
    10'b0010100101,
    10'b0100000001,
    10'b0101011001,
    10'b0101010101,
    10'b1000001001,
    10'b0001011110,
    10'b1000000111,
    10'b0001100100,
    10'b0111100100,
    10'b0011100100,
    10'b0101100000,
    10'b0110100100,
    10'b0100000000,
    10'b1001000100,
    10'b0010010000,
    10'b0100001100,
    10'b0011011100,
    10'b1001010100,
    10'b0101011100,
    10'b0001010100,
    10'b1000100100,
    10'b1000100000,
    10'b0111010100,
    10'b0000011001,
    10'b1001000001,
    10'b0001100001,
    10'b0000001101,
    10'b0001010001,
    10'b0000000101,
    10'b0010001001,
    10'b1000011001,
    10'b0101000101,
    10'b0111100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b0111100011,
    10'b0001011100,
    10'b0101000000,
    10'b0011011100,
    10'b0101011100,
    10'b0000011000,
    10'b0011100100,
    10'b1000001000,
    10'b0101010100,
    10'b0100010000,
    10'b0111010000,
    10'b1001010100,
    10'b0001001001,
    10'b1000100001,
    10'b0100010101,
    10'b0001100101,
    10'b0101001001,
    10'b0000001001,
    10'b0000100101,
    10'b1001000101,
    10'b0000010001,
    10'b0110100101,
    10'b0100001101,
    10'b0000100001,
    10'b0110000101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111000110,
    10'b0001011111,
    10'b0110001100,
    10'b0001001000,
    10'b0100010100,
    10'b0000001000,
    10'b1000001000,
    10'b0110010100,
    10'b0001001100,
    10'b0110000000,
    10'b0110011000,
    10'b0011011000,
    10'b0011001000,
    10'b0111010000,
    10'b0100000000,
    10'b0100100000,
    10'b1000000001,
    10'b0000011101,
    10'b0011010001,
    10'b0111010101,
    10'b0001100101,
    10'b0001010001,
    10'b0011011101,
    10'b1001011101,
    10'b0000000101,
    10'b0010100001,
    10'b0101100001,
    10'b1000100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001001110,
    10'b1000100011,
    10'b0101000100,
    10'b0011000000,
    10'b0011011100,
    10'b1000010000,
    10'b0000001000,
    10'b0110100100,
    10'b1001010000,
    10'b0010100000,
    10'b1000000100,
    10'b1001100100,
    10'b0101100100,
    10'b0001001001,
    10'b1000011101,
    10'b0010100101,
    10'b1000010101,
    10'b0101011101,
    10'b0010011101,
    10'b1001000101,
    10'b0001011001,
    10'b0101011001,
    10'b0110000101,
    10'b1001001101,
    10'b0000100001,
    10'b0011011001,
    10'b0010000101,
    10'b0100000101,
    10'b0101100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000011111,
    10'b0011100100,
    10'b0101000100,
    10'b1000010100,
    10'b0000010000,
    10'b0000010100,
    10'b0101010100,
    10'b0000000100,
    10'b0100010000,
    10'b1001010000,
    10'b0110011000,
    10'b0000000000,
    10'b0000001100,
    10'b0010011000,
    10'b0111100000,
    10'b0001000001,
    10'b1001011001,
    10'b0111000001,
    10'b0101010001,
    10'b0001011001,
    10'b0011001001,
    10'b0111001101,
    10'b0010010101,
    10'b0001011101,
    10'b0001100001,
    10'b0010001101,
    10'b0111011101,
    10'b0101100001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111001010,
    10'b0001100011,
    10'b0000001000,
    10'b0111100100,
    10'b0110001000,
    10'b0111011000,
    10'b1001010000,
    10'b0010010000,
    10'b1000001000,
    10'b0111000000,
    10'b0000010000,
    10'b0010000000,
    10'b0001011000,
    10'b0100001000,
    10'b0111001101,
    10'b0000100001,
    10'b0000000101,
    10'b0011010101,
    10'b0010011001,
    10'b0010000101,
    10'b0000011101,
    10'b1000000001,
    10'b0110011001,
    10'b0100011001,
    10'b0110010001,
    10'b1000010101,
    10'b0101011001,
    10'b0110000101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0110000110,
    10'b0001100011,
    10'b0001100100,
    10'b0010011100,
    10'b0100100100,
    10'b0111100100,
    10'b0110100000,
    10'b0001001000,
    10'b0001001100,
    10'b1000010100,
    10'b0100001100,
    10'b0011100000,
    10'b0010010000,
    10'b0100000100,
    10'b1000100100,
    10'b1001001100,
    10'b0000000100,
    10'b0110000000,
    10'b1001010000,
    10'b0110000001,
    10'b0010100001,
    10'b0001011001,
    10'b0101010001,
    10'b1000000001,
    10'b1000011101,
    10'b1001100101,
    10'b0000100101,
    10'b0100001001,
    10'b0101011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0111000110,
    10'b0010100011,
    10'b1001100100,
    10'b1000001000,
    10'b0001011100,
    10'b0100001100,
    10'b0101000000,
    10'b0111100100,
    10'b0001100100,
    10'b0111000000,
    10'b0111011000,
    10'b1001010100,
    10'b0110001001,
    10'b0011100101,
    10'b0000000001,
    10'b0111010101,
    10'b0100011101,
    10'b0101010101,
    10'b0110011001,
    10'b0010100101,
    10'b0010010101,
    10'b0100010101,
    10'b0101011001,
    10'b0100000101,
    10'b0100001001,
    10'b0111011101,
    10'b0000001001,
    10'b0011011101,
    10'b1001010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001110,
    10'b0001100011,
    10'b0110001100,
    10'b0010001000,
    10'b1001000100,
    10'b0011001100,
    10'b0111100000,
    10'b1001000000,
    10'b0001010000,
    10'b0101100000,
    10'b1001001000,
    10'b0111001001,
    10'b0000100001,
    10'b0101000001,
    10'b0100100001,
    10'b1001100001,
    10'b0000001001,
    10'b0100011001,
    10'b0111011101,
    10'b0010000001,
    10'b0010100001,
    10'b1001010001,
    10'b0100000101,
    10'b0101001001,
    10'b0010000101,
    10'b1001100101,
    10'b0001011001,
    10'b0100000001,
    10'b0101100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b1000011111,
    10'b0011011100,
    10'b1001100100,
    10'b0000100100,
    10'b1001011100,
    10'b0110000000,
    10'b1000000000,
    10'b0011000000,
    10'b0001000000,
    10'b0001001001,
    10'b0111100001,
    10'b0000001001,
    10'b0101001101,
    10'b0100010101,
    10'b0111000001,
    10'b0111000101,
    10'b0000010001,
    10'b1000001101,
    10'b1001100001,
    10'b1000010101,
    10'b0010100001,
    10'b0110011101,
    10'b0101011101,
    10'b0111001001,
    10'b0010010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0110001000,
    10'b0100000000,
    10'b0000000100,
    10'b0010100100,
    10'b0011100100,
    10'b0000011100,
    10'b0110010100,
    10'b1000010000,
    10'b0101000100,
    10'b0010000100,
    10'b0111100000,
    10'b0010011100,
    10'b1001001100,
    10'b0001100000,
    10'b0010001100,
    10'b1000001000,
    10'b0011001000,
    10'b0111011101,
    10'b0000001001,
    10'b0001011101,
    10'b0000010101,
    10'b0101100101,
    10'b0100000101,
    10'b0100001001,
    10'b0110011101,
    10'b0100010001,
    10'b1001000101,
    10'b1001000001,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001011011,
    10'b0110100100,
    10'b0000011100,
    10'b0001010000,
    10'b0011000100,
    10'b0001000000,
    10'b0111011100,
    10'b0101000100,
    10'b0001100000,
    10'b0110001000,
    10'b0100100000,
    10'b1000000001,
    10'b0001010101,
    10'b0001011101,
    10'b0101000001,
    10'b0000100001,
    10'b0010001001,
    10'b0011010001,
    10'b0100010101,
    10'b0111100101,
    10'b0110100001,
    10'b0011001101,
    10'b0000011001,
    10'b1001001101,
    10'b0001001101,
    10'b0000001101,
    10'b0101010101,
    10'b0110010001,
    10'b1001000001,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0011000111,
    10'b1000001100,
    10'b1000010000,
    10'b1000000100,
    10'b0010011000,
    10'b1001001100,
    10'b0001010000,
    10'b0111100100,
    10'b0111100000,
    10'b0101000000,
    10'b0010010000,
    10'b1000100100,
    10'b1000100101,
    10'b0100001001,
    10'b0110011001,
    10'b0000011101,
    10'b0110001001,
    10'b0000011001,
    10'b0001000101,
    10'b0100001101,
    10'b1001010101,
    10'b0010010101,
    10'b0111010101,
    10'b0000100101,
    10'b0111001101,
    10'b1001001001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001000110,
    10'b1000011011,
    10'b0100001000,
    10'b0110001000,
    10'b0100000000,
    10'b1001011100,
    10'b0010000000,
    10'b1000001100,
    10'b0000100000,
    10'b0100010100,
    10'b0000010000,
    10'b0000100100,
    10'b0000001001,
    10'b1001010101,
    10'b0101010101,
    10'b0111001001,
    10'b0001011101,
    10'b0000011101,
    10'b0011000101,
    10'b1000011101,
    10'b1001001001,
    10'b0111000001,
    10'b0001011001,
    10'b0100100001,
    10'b0001000001,
    10'b0111011001,
    10'b0001100001,
    10'b0011010101,
    10'b0101100101,
    10'b1000001001,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001111,
    10'b0000000000,
    10'b0011000000,
    10'b1001001100,
    10'b0001000100,
    10'b0000001000,
    10'b0111000100,
    10'b0010100000,
    10'b0000011000,
    10'b0100000000,
    10'b0010100100,
    10'b0100011100,
    10'b1000001000,
    10'b0101100100,
    10'b0111100001,
    10'b0010001001,
    10'b0110100101,
    10'b1000011001,
    10'b0110000001,
    10'b0101010101,
    10'b0100000101,
    10'b0001011101,
    10'b0111100101,
    10'b1000010101,
    10'b0010010101,
    10'b0111001101,
    10'b0101010001,
    10'b1000010001,
    10'b0001001001,
    10'b1111111100,
    10'b1111111100,
    10'b0001011110,
    10'b0111000111,
    10'b0100001000,
    10'b0111001100,
    10'b1000000000,
    10'b0101001000,
    10'b1001001000,
    10'b0000001000,
    10'b1001000100,
    10'b0111000000,
    10'b1000100100,
    10'b0111100000,
    10'b1001010100,
    10'b0011000100,
    10'b0100001100,
    10'b0011010100,
    10'b1000000100,
    10'b1001011100,
    10'b0000100001,
    10'b0111000001,
    10'b0011000001,
    10'b1001000001,
    10'b0110011001,
    10'b0001000101,
    10'b1000001001,
    10'b0100000001,
    10'b0001001001,
    10'b0000001101,
    10'b0000010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000100010,
    10'b0001001011,
    10'b0101010100,
    10'b0101000100,
    10'b1000001000,
    10'b1001011100,
    10'b0111011000,
    10'b0011011000,
    10'b0101011000,
    10'b0110011100,
    10'b0000000100,
    10'b1001001100,
    10'b0111000000,
    10'b0100100100,
    10'b1001011101,
    10'b0001001101,
    10'b0100011101,
    10'b0001011001,
    10'b1000010001,
    10'b0010100101,
    10'b0000011101,
    10'b0111010001,
    10'b1000000001,
    10'b0000010001,
    10'b0000011001,
    10'b0000100101,
    10'b0011001101,
    10'b0111001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001100011,
    10'b1001100000,
    10'b0000001000,
    10'b0100010100,
    10'b0111011000,
    10'b1001001000,
    10'b1001011000,
    10'b0010010000,
    10'b0110010100,
    10'b0111100100,
    10'b0100100100,
    10'b0101000100,
    10'b1000000101,
    10'b0010100001,
    10'b1001010001,
    10'b0101100101,
    10'b0110011101,
    10'b1001010101,
    10'b0111001101,
    10'b0100001101,
    10'b0101100001,
    10'b0011010101,
    10'b0110001001,
    10'b0010010101,
    10'b0110100001,
    10'b0000001101,
    10'b1000010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000000111,
    10'b0011100000,
    10'b0010010100,
    10'b0100100000,
    10'b0101100100,
    10'b0101010100,
    10'b0110010100,
    10'b0000011100,
    10'b0000010100,
    10'b0000001100,
    10'b0100000100,
    10'b0001000100,
    10'b1001100000,
    10'b0001100101,
    10'b0111000101,
    10'b0110001101,
    10'b0100100101,
    10'b0000000101,
    10'b0011010101,
    10'b0010011001,
    10'b0011100101,
    10'b1001010001,
    10'b1001011001,
    10'b0011000001,
    10'b1001010101,
    10'b0110100101,
    10'b0001000001,
    10'b0000010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0010100011,
    10'b0110000000,
    10'b0000001000,
    10'b0000010100,
    10'b1001100000,
    10'b0111001100,
    10'b0100010000,
    10'b0010010100,
    10'b0010001000,
    10'b0101000100,
    10'b0011010000,
    10'b0000011100,
    10'b0010100100,
    10'b1000011000,
    10'b0001011100,
    10'b0101010000,
    10'b0101010100,
    10'b0010011100,
    10'b0011010100,
    10'b1001000101,
    10'b0011100001,
    10'b1000000101,
    10'b0100100001,
    10'b0011001001,
    10'b1001011001,
    10'b1001001101,
    10'b0000000101,
    10'b0000001101,
    10'b0011100101,
    10'b0111011001,
    10'b0010000001,
    10'b1000001010,
    10'b0001100011,
    10'b0011000000,
    10'b0011011000,
    10'b0000011100,
    10'b0010011000,
    10'b0010001000,
    10'b0100000000,
    10'b1001011000,
    10'b1000100100,
    10'b0010001100,
    10'b0000001100,
    10'b0100010000,
    10'b1001010100,
    10'b0010000000,
    10'b0000100000,
    10'b0001011000,
    10'b0100100100,
    10'b1000001101,
    10'b0000011101,
    10'b1001001101,
    10'b0001001101,
    10'b0110100101,
    10'b0110100001,
    10'b1000010001,
    10'b0000010001,
    10'b0100011001,
    10'b0000000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b0111000111,
    10'b0001000000,
    10'b0110100000,
    10'b0100000100,
    10'b0101001000,
    10'b0101010100,
    10'b0000011000,
    10'b0111011000,
    10'b1000100000,
    10'b0110011000,
    10'b0001010000,
    10'b1000000000,
    10'b1001011000,
    10'b0000100101,
    10'b0110000001,
    10'b0011010001,
    10'b0100000001,
    10'b0101011101,
    10'b0111001001,
    10'b1000001101,
    10'b0011100001,
    10'b0001000101,
    10'b0110000101,
    10'b0100010101,
    10'b0010001101,
    10'b0101100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000011111,
    10'b0101001000,
    10'b0011100000,
    10'b0111001100,
    10'b0011000000,
    10'b0101100100,
    10'b0100100000,
    10'b0000100000,
    10'b0110000100,
    10'b1001100100,
    10'b0011000001,
    10'b0111011001,
    10'b0010100101,
    10'b0011011001,
    10'b0010100001,
    10'b1000000101,
    10'b0011000101,
    10'b0101011001,
    10'b0110100001,
    10'b0101001101,
    10'b0110010101,
    10'b0001001001,
    10'b0001000001,
    10'b0100001101,
    10'b0010011101,
    10'b0100000001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010100010,
    10'b0111000111,
    10'b1000011000,
    10'b0101010100,
    10'b1001011100,
    10'b1000000000,
    10'b0011100000,
    10'b0011000100,
    10'b0110011100,
    10'b0000000100,
    10'b0100000000,
    10'b0001000000,
    10'b1001010100,
    10'b0111000000,
    10'b0011001100,
    10'b0000010000,
    10'b0111100100,
    10'b1001010000,
    10'b0110010000,
    10'b0111011000,
    10'b0011011101,
    10'b1000001001,
    10'b0100100101,
    10'b0101010001,
    10'b0110000001,
    10'b0100011001,
    10'b0010000001,
    10'b0001011001,
    10'b0011011001,
    10'b0101100101,
    10'b0110001101,
    10'b1111111100,
    10'b0001001010,
    10'b1000011111,
    10'b1000010100,
    10'b0100000000,
    10'b0110011000,
    10'b0100010100,
    10'b0000000000,
    10'b0110011100,
    10'b0010010000,
    10'b0010011000,
    10'b0101011100,
    10'b0110100100,
    10'b0101100100,
    10'b0100011000,
    10'b0010000101,
    10'b0111100001,
    10'b0000100101,
    10'b1000001001,
    10'b0010010101,
    10'b0011001101,
    10'b0110100001,
    10'b1001001001,
    10'b0110010001,
    10'b0111001101,
    10'b1001011101,
    10'b0001011101,
    10'b0011100001,
    10'b0011011001,
    10'b1000001101,
    10'b0101001001,
    10'b0111011101,
    10'b1111111100,
    10'b0001000110,
    10'b1000100011,
    10'b0101001000,
    10'b0111000100,
    10'b0111100100,
    10'b0011010100,
    10'b0011001000,
    10'b0100001000,
    10'b0000010100,
    10'b0110011100,
    10'b0010010100,
    10'b0110000000,
    10'b0000000001,
    10'b0111011101,
    10'b0100011001,
    10'b0010011101,
    10'b0100100101,
    10'b0010011001,
    10'b0000001001,
    10'b1000011001,
    10'b1001000001,
    10'b0111100001,
    10'b0001100101,
    10'b1000010101,
    10'b0110001001,
    10'b0111010101,
    10'b1001001001,
    10'b0010100001,
    10'b0011010001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0010000110,
    10'b1000100011,
    10'b1001100000,
    10'b0011100100,
    10'b0011001000,
    10'b0100001100,
    10'b0010010100,
    10'b0100100100,
    10'b0011011100,
    10'b0001100100,
    10'b0110010100,
    10'b0111011000,
    10'b0111001000,
    10'b0010010000,
    10'b0111011100,
    10'b1000100100,
    10'b0010001001,
    10'b1001100001,
    10'b0101010101,
    10'b0110100101,
    10'b0010100001,
    10'b1000000101,
    10'b1000010001,
    10'b1001010001,
    10'b0000011001,
    10'b0101001101,
    10'b0001001101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001011111,
    10'b1000000000,
    10'b0110000100,
    10'b1001010100,
    10'b0110011100,
    10'b0110000000,
    10'b0001000000,
    10'b1000011100,
    10'b0011011100,
    10'b0000000000,
    10'b1000000001,
    10'b0010011001,
    10'b0100011101,
    10'b0011011001,
    10'b0110011001,
    10'b1000100001,
    10'b0100011001,
    10'b0100001001,
    10'b0000011001,
    10'b0111011001,
    10'b0110010101,
    10'b0000100101,
    10'b0010000101,
    10'b0010100101,
    10'b0101011101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0011100011,
    10'b0101100100,
    10'b1001010000,
    10'b0000100100,
    10'b0001000000,
    10'b0010010000,
    10'b0010100100,
    10'b0010010100,
    10'b0110100000,
    10'b1001000000,
    10'b0001011100,
    10'b1001001001,
    10'b0100100001,
    10'b0011000001,
    10'b1000010101,
    10'b0001000101,
    10'b0111001001,
    10'b1000010001,
    10'b1001100101,
    10'b0111011001,
    10'b1000001101,
    10'b0001010101,
    10'b0001100101,
    10'b0010011001,
    10'b0000000101,
    10'b0111001101,
    10'b1000000001,
    10'b0000000001,
    10'b0110010101,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b1000001111,
    10'b0011001000,
    10'b0101011100,
    10'b0001100100,
    10'b0001010000,
    10'b0111010100,
    10'b0000010100,
    10'b0110000100,
    10'b0100001100,
    10'b0000100100,
    10'b0000011000,
    10'b0011001100,
    10'b1001100100,
    10'b1000010100,
    10'b0011100000,
    10'b0100011100,
    10'b1000011000,
    10'b0110000000,
    10'b0010100001,
    10'b1000001001,
    10'b0010000001,
    10'b0001011001,
    10'b0000010001,
    10'b0011011101,
    10'b0110001101,
    10'b0110100101,
    10'b1001010001,
    10'b0111011101,
    10'b0111001001,
    10'b0010011101,
    10'b0100100001,
    10'b0110000110,
    10'b0001100011,
    10'b0100011000,
    10'b0000011000,
    10'b1001001000,
    10'b0011001000,
    10'b0001100100,
    10'b1000000100,
    10'b1000001100,
    10'b0111011000,
    10'b0000000100,
    10'b0111000001,
    10'b0000100001,
    10'b1001100101,
    10'b1001010101,
    10'b0101000101,
    10'b0000010101,
    10'b0000011101,
    10'b0000010001,
    10'b0110010001,
    10'b0111001101,
    10'b0100001101,
    10'b0010100001,
    10'b1000011101,
    10'b0111011101,
    10'b0011000101,
    10'b0101011101,
    10'b0010011001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0001100011,
    10'b0110010100,
    10'b0100100100,
    10'b1000011100,
    10'b0100000100,
    10'b0100010000,
    10'b0110000000,
    10'b0111011100,
    10'b0011011000,
    10'b0110010000,
    10'b0010000100,
    10'b0011000100,
    10'b1001000000,
    10'b1001011100,
    10'b0000010000,
    10'b1001000100,
    10'b0111001000,
    10'b1000100000,
    10'b1001000001,
    10'b0001100101,
    10'b0111100001,
    10'b0001001001,
    10'b0100001001,
    10'b0010100101,
    10'b0101000101,
    10'b0000011101,
    10'b1001010101,
    10'b1001001101,
    10'b0000010101,
    10'b1111111100,
    10'b1111111100,
    10'b0001100010,
    10'b0110000111,
    10'b1000001100,
    10'b0110010100,
    10'b0001011100,
    10'b0011011000,
    10'b0101011000,
    10'b0011011100,
    10'b0101010100,
    10'b1001010100,
    10'b1001100000,
    10'b0010011101,
    10'b0101000001,
    10'b0111000101,
    10'b1000011101,
    10'b1000010101,
    10'b0101010001,
    10'b0011100101,
    10'b0111010101,
    10'b0000010101,
    10'b0101001101,
    10'b0100100001,
    10'b0101011101,
    10'b0101000101,
    10'b0100000001,
    10'b0000100101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1000000110,
    10'b0011100011,
    10'b0011001000,
    10'b0010100100,
    10'b0001000000,
    10'b0011011100,
    10'b0111010100,
    10'b0101001000,
    10'b0110001100,
    10'b0100001000,
    10'b1001001000,
    10'b0101000100,
    10'b0110100100,
    10'b0000001100,
    10'b1001010100,
    10'b0011000100,
    10'b1001011100,
    10'b1000100000,
    10'b0000011100,
    10'b0001011000,
    10'b1001000101,
    10'b0010011101,
    10'b0111001101,
    10'b0111001001,
    10'b0000000101,
    10'b0110100001,
    10'b0111010001,
    10'b0000010101,
    10'b1001100001,
    10'b1000010001,
    10'b0101100101,
    10'b0000100001,
    10'b0001011110,
    10'b0111000111,
    10'b0011001100,
    10'b1000000100,
    10'b0110100000,
    10'b1000011000,
    10'b0100011100,
    10'b0101010000,
    10'b1001010100,
    10'b0000010000,
    10'b1000100100,
    10'b1001100100,
    10'b0000011000,
    10'b0100010100,
    10'b0010000000,
    10'b0000100100,
    10'b0100100100,
    10'b0011011100,
    10'b0010100001,
    10'b0110000101,
    10'b0110011001,
    10'b0010011101,
    10'b1001000101,
    10'b0011011001,
    10'b1000001001,
    10'b1001001101,
    10'b0000000101,
    10'b0101010101,
    10'b0000000001,
    10'b1000010101,
    10'b1111111100,
    10'b1111111100,
    10'b1000001010,
    10'b0001100011,
    10'b0100010000,
    10'b0010000000,
    10'b0111010100,
    10'b1001000100,
    10'b0110010000,
    10'b1000010000,
    10'b0100000100,
    10'b0100001100,
    10'b0110001000,
    10'b0001000100,
    10'b0010010100,
    10'b0100000000,
    10'b1001000101,
    10'b0000100101,
    10'b0111001001,
    10'b0001011001,
    10'b0011100001,
    10'b0111011101,
    10'b1001100001,
    10'b0100010101,
    10'b1000001101,
    10'b0011001001,
    10'b0111000101,
    10'b0110000101,
    10'b0000100001,
    10'b0001001001,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b0110000110,
    10'b0001100011,
    10'b0101010000,
    10'b0111011100,
    10'b1000000000,
    10'b0111010000,
    10'b1000010100,
    10'b1000100100,
    10'b0001010000,
    10'b0001011100,
    10'b0101100000,
    10'b0010010100,
    10'b0010010000,
    10'b0100001000,
    10'b0111001001,
    10'b0000100001,
    10'b0001000101,
    10'b0010100101,
    10'b1001010101,
    10'b0101001001,
    10'b0011011001,
    10'b0101000101,
    10'b0111100001,
    10'b0000000101,
    10'b0010011101,
    10'b0100010101,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
    10'b1111111100,
};

endmodule
